module transmission_gate(inout a, inout b, input c);
   tranif1(a, b, c);
endmodule
